`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.12.2023 14:32:56
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(
    input clkvga, clk,
    //input [7:0] entera, enterd,
    input [15:0] enter,
    input clk2,clk3,          // 100MHz on Basys 3
    input reset,rst,        // btnC on Basys 3
    output hsync,       // to VGA connector
    output vsync,       // to VGA connector
    output [11:0] rgb   // to DAC, to VGA connector
    );
    
    // signals
    wire [9:0] w_x, w_y;
    wire w_video_on, w_p_tick;
    reg [11:0] rgb_reg;
    wire [11:0] rgb_next;
    
    // VGA Controller
    vga_controller vga(.clk_100MHz(clkvga), .reset(reset), .hsync(hsync), .vsync(vsync),
                       .video_on(w_video_on), .p_tick(w_p_tick), .x(w_x), .y(w_y));
    // Text Generation Circuit
    //ascii_test at(.clkvga(clkvga), .entera(entera), .enterd(enterd), .clk2(clk2), .clk(clk),  .video_on(w_video_on), .x(w_x), .y(w_y), .rgb(rgb_next) );
    ascii_test at(.clkvga(clkvga), .enter(enter), .rst(rst), .clk2(clk2), .clk3(clk3), .clk(clk), .video_on(w_video_on), .x(w_x), .y(w_y), .rgb(rgb_next) );
    //ascii_test at(.clkvga(clkvga), .enter(enter), .rst(rst),.clk2(clk2), .clk3(clk3),  .video_on(w_video_on), .x(w_x), .y(w_y), .rgb(rgb_next) );
    
    // rgb buffer
    always @(posedge clkvga)
        if(w_p_tick)
            rgb_reg <= rgb_next;
            
    // output
    assign rgb = rgb_reg;
      
endmodule